library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package global_configuration is
  
  constant c_FPGA_MANUFACTURER : STRING  := "GOWIN";
  constant c_CLOCK_FREQUENCY   : natural := 48000000;
  
end package global_configuration;
 
package body global_configuration is
 
end package body global_configuration;